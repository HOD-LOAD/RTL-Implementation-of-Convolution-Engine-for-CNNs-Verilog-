module hello;
  initial begin
    $display("Hello, Icarus Verilog is working!");
    $finish;
  end
endmodule
